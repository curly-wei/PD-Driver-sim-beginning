.title Equivalent photodiode model

	.subckt PDMod IpdN IpdP kCpd=11pF kRpd=38G
		******
		** kIpd: Equivalent current source of photodiode /Constant
		** kCpd: Equivalent capacitor of photodiode /Constant
		** kRs: Equivalent Resistor of photodiode /Constant
		** IpdP: Photodiode current output, N-type (Cathod)
		** IpdN: Photodiode current output, P-type (Anode)
		******	
		
		C_pd IpdP IpdN {kCpd}
		R_pd IpdP IpdN {kRpd}
		
		******
		** Pulse for emulate PD current output
		** pulse( V_init V_pulse T_delay T_risetime T_falltime PulseWidth Period )
		I_pd IpdN IpdP pulse( 0 10nA 0ns 20ns 20ns 40ns 300us )
		******
	
	.ends
.end
