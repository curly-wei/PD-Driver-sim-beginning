.title I/V Converter for PD-Driver

  .include lib/OPAx192/OPAx192.LIB
  .subckt IVCvT_OPA192 Ii Vo Vdd Vss kCfb=2.7pF kRfb=1Meg kRbu=42k kRbd=3k
		******	
		** Implement IV converter with OPA192
		** kCpd: Equivelated capacitor of photodiode /Constant 
		** kCfb: Feedback capacitor /Constant 
		** kRfb: Feedback resistor /Constant 
		** kRbu: Bias resistor(up) for voltage divider numerator /Constant 
		** kRbd: Bias resistor(down) for voltage divider denominator /Constant 
		** Ii: Current source input 
		** Vo: Volatge output 
		** Vcc: System power high
		** Vss: System power low 	
		****** 
		C_fb Ii Vo {kCfb}
		R_fb Ii Vo {kRfb}
		R_bu Vdd nVbias {kRbu}
		R_bd nVbias Vss {kRbd}
		X_OPA192 nVbias Ii Vdd Vss Vo OPAx192
  .ends

	.include lib/OPA810/opa810_a.lib
  .subckt IVCvT_OPA810 Ii Vo Vdd Vss kCfb=2.7pF kRfb=1Meg kRbu=42k kRbd=3k
		******	
		** Implement IV converter with OPA810
		** kCpd: Equivelated capacitor of photodiode /Constant 
		** kCfb: Feedback capacitor /Constant 
		** kRfb: Feedback resistor /Constant 
		** kRbu: Bias resistor(up) for voltage divider numerator /Constant 
		** kRbd: Bias resistor(down) for voltage divider denominator /Constant 
		** Ii: Current source input 
		** Vo: Volatge output 
		** Vcc: System power high
		** Vss: System power low 	
		******
		C_fb Ii Vo {kCfb}
		R_fb Ii Vo {kRfb}
		R_bu Vdd nVbias {kRbu}
		R_bd nVbias Vss {kRbd}
		X_OPA810 nVbias Ii Vo Vdd Vss OPA810
  .ends

	.include lib/LMH6601/LMH6601.MOD
  .subckt IVCvT_LMH6601 Ii Vo Vdd Vss kCfb=2.7pF kRfb=1Meg kRbu=42k kRbd=3k
		******	
		** Implement IV converter with LMH6601
		** kCpd: Equivelated capacitor of photodiode /Constant 
		** kCfb: Feedback capacitor /Constant 
		** kRfb: Feedback resistor /Constant 
		** kRbu: Bias resistor(up) for voltage divider numerator /Constant 
		** kRbd: Bias resistor(down) for voltage divider denominator /Constant 
		** Ii: Current source input 
		** Vo: Volatge output 
		** Vcc: System power high
		** Vss: System power low 	
		******
		C_fb Ii Vo {kCfb}
		R_fb Ii Vo {kRfb}
		R_bu Vdd nVbias {kRbu}
		R_bd nVbias Vss {kRbd}
		X_LMH6601 nVbias Ii Vdd Vss Vo LMH6601
  .ends
	
	.include lib/ada4817/ada4817.cir
  .subckt IVCvT_ADA4817 Ii Vo Vdd Vss kCfb=27pF kRfb=1Meg kRbu=42k kRbd=3k
		******	
		** Implement IV converter with ADA4817
		** kCpd: Equivelated capacitor of photodiode /Constant 
		** kCfb: Feedback capacitor /Constant 
		** kRfb: Feedback resistor /Constant 
		** kRbu: Bias resistor(up) for voltage divider numerator /Constant 
		** kRbd: Bias resistor(down) for voltage divider denominator /Constant 
		** Ii: Current source input 
		** Vo: Volatge output 
		** Vcc: System power high
		** Vss: System power low 	
		****** 
		C_fb Ii Vfb {kCfb}  
		R_fb Ii Vfb {kRfb}
		R_bu Vdd nVbias {kRbu}
		R_bd nVbias Vss {kRbd} 
		X_ADA4817 nVbias Ii Vdd Vss Vo Vfb Vdd ADA4817
  .ends


.end
