.title Testbench for PD-Driver
  .include IVCvT_OPA810.cir
  .include PDMod.cir

  VCC 5v0 GND DC 5V
  
  X_IVCvT nPD_Io nIVCvt_Vo 5v0 GND IVCvT_OPA810 kCfb=20pF kRfb=1k
  X_PDMod nPD_Io GND PDMod
  
  .control
    * set ctrl var
    set tran_data_out_filename="pd-tran-opa810.ssv"
    * Transient Analyze
    tran 5n 5u ;tran <step> <stop>
    * Save data to ssv file
    wrdata $tran_data_out_filename V(nIVCvt_Vo) 
    ssd
    exit
  .endc



.end
