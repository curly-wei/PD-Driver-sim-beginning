.title Equivalent photodiode model

	.subckt pd_model IpdCathod IpdAnode kCpd=400pF kRpd=38G
		******
		** kIpd: Equivalent current source of photodiode /Constant
		** kCpd: Equivalent capacitor of photodiode /Constant
		** kRs: Equivalent Resistor of photodiode /Constant
		** IpdCathod: Photodiode current output, Cathod
		** IpdAnode: Photodiode current output, Anode
		******	
		
		C_pd IpdCathod IpdAnode {kCpd}
		R_pd IpdCathod IpdAnode {kRpd}
		
		******
		** Pulse for emulate PD current output
		** pulse( V_init V_pulse T_delay T_risetime T_falltime PulseWidth Period )
		I_pd IpdCathod IpdAnode pulse( 0 1uA 100ns 6us 6us 10us 3000us )
		******
	
	.ends
.end
