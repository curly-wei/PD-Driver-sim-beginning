.title Testbench for PD-Driver
  .include IVCvT_ADA4817.cir
  .include PDMod.cir

 
  VCC 5V0 GND DC 5V

  X_IVCvT nPD_Io nIVCvt_Vo 5V0 GND IVCvT_ADA4817 kCfb=0 kRfb=1Meg
  X_PDMod nPD_Io GND PDMod
   
 
  .control
    * set ctrl var
    set tran_data_out_filename="pd-tran-ada4817.ssv"
    * Transient Analyze
    tran 1n 10u ;tran <step> <stop>
    listing
    * plot V(nIVCvt_Vo) 
    * Save data to ssv file
    wrdata $tran_data_out_filename V(nIVCvt_Vo) 
    exit
  .endc



.end
