** Profile: "SCHEMATIC1-ac_sweep"  [ C:\Users\a0232073\Desktop\GWL_Models\OPA810\AppendScript\opa810_pspice\opa810_pspice-pspicefiles\schematic1\ac_sweep.sim ] 

** Creating circuit file "ac_sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../opa810_a.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpiceTIPSpice_Install\17.4.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 1n 
.OPTIONS ADVCONV
.PROBE64 N([OUT])
.PROBE64 N([IN+])
.INC "..\SCHEMATIC1.net" 


.END
