.title Testbench for PD-Driver
  .include ../IVCvT.cir
  .include ../PDMod.cir


  VCC 4v5 GND DC 4.5V
  
  X_IVCvT nPD_Io nIVCvt_Vo 4v5 GND IVCvT_OPA355 kCfb=100fF kRfb=100Meg
  X_PDMod nPD_Io GND PDMod
  

  .control
    * set ctrl var
    set tran_data_out_filename="pd-tran-opa355.ssv"
    * Transient Analyze
    tran 5n 50u ;tran <step> <stop>
    * Save data to ssv file 
    wrdata $tran_data_out_filename V(nIVCvt_Vo) 
    exit
  .endc



.end
