.title impl_OPAx192_cir
  .include OPAx192/OPAx192.LIB
  .subckt impl_OPAx192_cir Ii Vo Vdd Vss kCfb=2.7pF kRfb=1Meg kRbu=4k kRbd=1k
		******	
		** kCpd: Equivelated capacitor of photodiode /Constant 
		** kCfb: Feedback capacitor /Constant 
		** kRfb: Feedback resistor /Constant 
		** kRbu: Bias resistor(up) for voltage divider numerator /Constant 
		** kRbd: Bias resistor(down) for voltage divider denominator /Constant 
		** Ii: Current source input 
		** Vo: Volatge output 
		** Vcc: System power high
		** Vss: System power low 	
		******
		C_fb Ii Vo {kCfb}
		R_fb Ii Vo {kRfb}
		R_bu Vdd n_bias {kRbu}
		R_bd n_bias Vss {kRbd}
		X_OPA192 n_bias Ii Vdd Vss Vo OPAx192
  .ends

.end
