.title I/V Converter for PD-Driver
  .include lib/LMH6601/LMH6601.MOD
  .subckt IVCvT_LMH6601 Ii Vo Vdd Vss kCfb=2.7pF kRfb=1Meg kRbu=47k kRbd=3k
		******	
		** kCpd: Equivelated capacitor of photodiode /Constant 
		** kCfb: Feedback capacitor /Constant 
		** kRfb: Feedback resistor /Constant 
		** kRbu: Bias resistor(up) for voltage divider numerator /Constant 
		** kRbd: Bias resistor(down) for voltage divider denominator /Constant 
		** Ii: Current source input 
		** Vo: Volatge output 
		** Vcc: System power high
		** Vss: System power low 	
		******
		C_fb Ii Vo {kCfb}
		R_fb Ii Vo {kRfb}
		R_bu Vdd nVbias {kRbu}
		R_bd nVbias Vss {kRbd}
		X_LMH6601 nVbias Ii Vdd Vss Vo LMH6601
  .ends

.end
