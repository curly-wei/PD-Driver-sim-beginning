.title Testbench for OPAx192_cir
  .include impl_OPAx192_cir.cir
  .include pd_model.cir

  VCC 5v0 GND DC 5V

  X_opa192 n_pd_o n_Vout 5v0 GND impl_OPAx192_cir
  X_pd_model n_pd_o GND pd_model

  
	.control
  	tran 100n 200u
    run
    plot V(n_Vout) 
  .endc

.end
