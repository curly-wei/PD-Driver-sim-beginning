.title I/V Converter for PD-Driver
  .include lib/ada4817/ada4817.cir
  .subckt IVCvT_ADA4817 Ii Vo Vdd Vss kCfb=27pF kRfb=1Meg kRbu=47k kRbd=3k
		******	
		** kCpd: Equivelated capacitor of photodiode /Constant 
		** kCfb: Feedback capacitor /Constant 
		** kRfb: Feedback resistor /Constant 
		** kRbu: Bias resistor(up) for voltage divider numerator /Constant 
		** kRbd: Bias resistor(down) for voltage divider denominator /Constant 
		** Ii: Current source input 
		** Vo: Volatge output 
		** Vcc: System power high
		** Vss: System power low 	
		****** 
		C_fb Ii Vfb {kCfb}  
		R_fb Ii Vfb {kRfb}
		R_bu Vdd nVbias {kRbu}
		R_bd nVbias Vss {kRbd} 
		X_ADA4817 nVbias Ii Vdd Vss Vo Vfb Vdd ADA4817
  .ends

.end
