.title Testbench for PD-Driver
  .include IVCvT.cir
  .include PDMod.cir

  VCC 5v0 GND DC 5V

  X_IVCvT nPD_Io nIVCvt_Vo 5v0 GND IVCvT
  X_PDMod nPD_Io GND PDMod
  
  .control
    * set ctrl var
    set tran_data_out_filename="pd-tran.ssv"
    * Transient Analyze
    tran 0.1u 200u ;tran <step> <stop>
    * Save data to ssv file
    wrdata $tran_data_out_filename V(nIVCvt_Vo) 
    ssd
    exit
  .endc



.end
